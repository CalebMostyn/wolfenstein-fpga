module raycast(
	input wire [9:0]x_pixel, 	// currently drawn pixel x
	input wire [9:0]y_pixel, 	// currently drawn pixel y
	output wire [639:0]is_in_rays,
	output wire [1279:0]ray_colors
);

parameter BLACK = 2'd0,
			RED = 2'd1,
			GREEN = 2'd2,
			BLUE = 2'd3;

parameter MAX_HEIGHT = 480 - 200;

// Square: (x top left, y top left, width, height, x_pixel, y_pixel, is_in_rays[i])
square ray_0(0,100 + ((MAX_HEIGHT - 172) / 2),1,172, x_pixel, y_pixel, is_in_rays[0]);
assign ray_colors[1:0] = RED;
square ray_1(1,100 + ((MAX_HEIGHT - 172) / 2),1,172, x_pixel, y_pixel, is_in_rays[1]);
assign ray_colors[3:2] = RED;
square ray_2(2,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[2]);
assign ray_colors[5:4] = RED;
square ray_3(3,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[3]);
assign ray_colors[7:6] = RED;
square ray_4(4,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[4]);
assign ray_colors[9:8] = RED;
square ray_5(5,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[5]);
assign ray_colors[11:10] = RED;
square ray_6(6,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[6]);
assign ray_colors[13:12] = RED;
square ray_7(7,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[7]);
assign ray_colors[15:14] = RED;
square ray_8(8,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[8]);
assign ray_colors[17:16] = RED;
square ray_9(9,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[9]);
assign ray_colors[19:18] = RED;
square ray_10(10,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[10]);
assign ray_colors[21:20] = RED;
square ray_11(11,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[11]);
assign ray_colors[23:22] = RED;
square ray_12(12,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[12]);
assign ray_colors[25:24] = RED;
square ray_13(13,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[13]);
assign ray_colors[27:26] = RED;
square ray_14(14,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[14]);
assign ray_colors[29:28] = RED;
square ray_15(15,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[15]);
assign ray_colors[31:30] = RED;
square ray_16(16,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[16]);
assign ray_colors[33:32] = RED;
square ray_17(17,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[17]);
assign ray_colors[35:34] = RED;
square ray_18(18,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[18]);
assign ray_colors[37:36] = RED;
square ray_19(19,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[19]);
assign ray_colors[39:38] = RED;
square ray_20(20,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[20]);
assign ray_colors[41:40] = RED;
square ray_21(21,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[21]);
assign ray_colors[43:42] = RED;
square ray_22(22,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[22]);
assign ray_colors[45:44] = RED;
square ray_23(23,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[23]);
assign ray_colors[47:46] = RED;
square ray_24(24,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[24]);
assign ray_colors[49:48] = RED;
square ray_25(25,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[25]);
assign ray_colors[51:50] = RED;
square ray_26(26,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[26]);
assign ray_colors[53:52] = RED;
square ray_27(27,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[27]);
assign ray_colors[55:54] = RED;
square ray_28(28,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[28]);
assign ray_colors[57:56] = RED;
square ray_29(29,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[29]);
assign ray_colors[59:58] = RED;
square ray_30(30,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[30]);
assign ray_colors[61:60] = RED;
square ray_31(31,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[31]);
assign ray_colors[63:62] = RED;
square ray_32(32,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[32]);
assign ray_colors[65:64] = RED;
square ray_33(33,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[33]);
assign ray_colors[67:66] = RED;
square ray_34(34,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[34]);
assign ray_colors[69:68] = RED;
square ray_35(35,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[35]);
assign ray_colors[71:70] = RED;
square ray_36(36,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[36]);
assign ray_colors[73:72] = RED;
square ray_37(37,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[37]);
assign ray_colors[75:74] = RED;
square ray_38(38,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[38]);
assign ray_colors[77:76] = RED;
square ray_39(39,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[39]);
assign ray_colors[79:78] = RED;
square ray_40(40,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[40]);
assign ray_colors[81:80] = RED;
square ray_41(41,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[41]);
assign ray_colors[83:82] = RED;
square ray_42(42,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[42]);
assign ray_colors[85:84] = RED;
square ray_43(43,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[43]);
assign ray_colors[87:86] = RED;
square ray_44(44,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[44]);
assign ray_colors[89:88] = RED;
square ray_45(45,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[45]);
assign ray_colors[91:90] = RED;
square ray_46(46,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[46]);
assign ray_colors[93:92] = RED;
square ray_47(47,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[47]);
assign ray_colors[95:94] = RED;
square ray_48(48,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[48]);
assign ray_colors[97:96] = RED;
square ray_49(49,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[49]);
assign ray_colors[99:98] = RED;
square ray_50(50,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[50]);
assign ray_colors[101:100] = RED;
square ray_51(51,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[51]);
assign ray_colors[103:102] = RED;
square ray_52(52,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[52]);
assign ray_colors[105:104] = RED;
square ray_53(53,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[53]);
assign ray_colors[107:106] = RED;
square ray_54(54,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[54]);
assign ray_colors[109:108] = RED;
square ray_55(55,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[55]);
assign ray_colors[111:110] = RED;
square ray_56(56,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[56]);
assign ray_colors[113:112] = RED;
square ray_57(57,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[57]);
assign ray_colors[115:114] = RED;
square ray_58(58,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[58]);
assign ray_colors[117:116] = RED;
square ray_59(59,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[59]);
assign ray_colors[119:118] = RED;
square ray_60(60,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[60]);
assign ray_colors[121:120] = RED;
square ray_61(61,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[61]);
assign ray_colors[123:122] = RED;
square ray_62(62,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[62]);
assign ray_colors[125:124] = RED;
square ray_63(63,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[63]);
assign ray_colors[127:126] = RED;
square ray_64(64,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[64]);
assign ray_colors[129:128] = RED;
square ray_65(65,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[65]);
assign ray_colors[131:130] = RED;
square ray_66(66,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[66]);
assign ray_colors[133:132] = RED;
square ray_67(67,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[67]);
assign ray_colors[135:134] = RED;
square ray_68(68,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[68]);
assign ray_colors[137:136] = RED;
square ray_69(69,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[69]);
assign ray_colors[139:138] = RED;
square ray_70(70,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[70]);
assign ray_colors[141:140] = RED;
square ray_71(71,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[71]);
assign ray_colors[143:142] = RED;
square ray_72(72,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[72]);
assign ray_colors[145:144] = RED;
square ray_73(73,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[73]);
assign ray_colors[147:146] = RED;
square ray_74(74,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[74]);
assign ray_colors[149:148] = RED;
square ray_75(75,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[75]);
assign ray_colors[151:150] = RED;
square ray_76(76,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[76]);
assign ray_colors[153:152] = RED;
square ray_77(77,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[77]);
assign ray_colors[155:154] = RED;
square ray_78(78,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[78]);
assign ray_colors[157:156] = RED;
square ray_79(79,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[79]);
assign ray_colors[159:158] = RED;
square ray_80(80,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[80]);
assign ray_colors[161:160] = RED;
square ray_81(81,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[81]);
assign ray_colors[163:162] = RED;
square ray_82(82,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[82]);
assign ray_colors[165:164] = RED;
square ray_83(83,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[83]);
assign ray_colors[167:166] = RED;
square ray_84(84,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[84]);
assign ray_colors[169:168] = RED;
square ray_85(85,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[85]);
assign ray_colors[171:170] = RED;
square ray_86(86,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[86]);
assign ray_colors[173:172] = RED;
square ray_87(87,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[87]);
assign ray_colors[175:174] = RED;
square ray_88(88,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[88]);
assign ray_colors[177:176] = RED;
square ray_89(89,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[89]);
assign ray_colors[179:178] = RED;
square ray_90(90,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[90]);
assign ray_colors[181:180] = RED;
square ray_91(91,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[91]);
assign ray_colors[183:182] = RED;
square ray_92(92,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[92]);
assign ray_colors[185:184] = RED;
square ray_93(93,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[93]);
assign ray_colors[187:186] = RED;
square ray_94(94,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[94]);
assign ray_colors[189:188] = RED;
square ray_95(95,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[95]);
assign ray_colors[191:190] = RED;
square ray_96(96,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[96]);
assign ray_colors[193:192] = RED;
square ray_97(97,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[97]);
assign ray_colors[195:194] = RED;
square ray_98(98,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[98]);
assign ray_colors[197:196] = RED;
square ray_99(99,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[99]);
assign ray_colors[199:198] = RED;
square ray_100(100,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[100]);
assign ray_colors[201:200] = RED;
square ray_101(101,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[101]);
assign ray_colors[203:202] = RED;
square ray_102(102,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[102]);
assign ray_colors[205:204] = RED;
square ray_103(103,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[103]);
assign ray_colors[207:206] = RED;
square ray_104(104,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[104]);
assign ray_colors[209:208] = RED;
square ray_105(105,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[105]);
assign ray_colors[211:210] = RED;
square ray_106(106,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[106]);
assign ray_colors[213:212] = RED;
square ray_107(107,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[107]);
assign ray_colors[215:214] = RED;
square ray_108(108,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[108]);
assign ray_colors[217:216] = RED;
square ray_109(109,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[109]);
assign ray_colors[219:218] = RED;
square ray_110(110,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[110]);
assign ray_colors[221:220] = RED;
square ray_111(111,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[111]);
assign ray_colors[223:222] = RED;
square ray_112(112,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[112]);
assign ray_colors[225:224] = RED;
square ray_113(113,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[113]);
assign ray_colors[227:226] = RED;
square ray_114(114,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[114]);
assign ray_colors[229:228] = RED;
square ray_115(115,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[115]);
assign ray_colors[231:230] = RED;
square ray_116(116,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[116]);
assign ray_colors[233:232] = RED;
square ray_117(117,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[117]);
assign ray_colors[235:234] = RED;
square ray_118(118,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[118]);
assign ray_colors[237:236] = RED;
square ray_119(119,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[119]);
assign ray_colors[239:238] = RED;
square ray_120(120,100 + ((MAX_HEIGHT - 172) / 2),1,172, x_pixel, y_pixel, is_in_rays[120]);
assign ray_colors[241:240] = RED;
square ray_121(121,100 + ((MAX_HEIGHT - 171) / 2),1,171, x_pixel, y_pixel, is_in_rays[121]);
assign ray_colors[243:242] = RED;
square ray_122(122,100 + ((MAX_HEIGHT - 170) / 2),1,170, x_pixel, y_pixel, is_in_rays[122]);
assign ray_colors[245:244] = RED;
square ray_123(123,100 + ((MAX_HEIGHT - 170) / 2),1,170, x_pixel, y_pixel, is_in_rays[123]);
assign ray_colors[247:246] = RED;
square ray_124(124,100 + ((MAX_HEIGHT - 169) / 2),1,169, x_pixel, y_pixel, is_in_rays[124]);
assign ray_colors[249:248] = RED;
square ray_125(125,100 + ((MAX_HEIGHT - 168) / 2),1,168, x_pixel, y_pixel, is_in_rays[125]);
assign ray_colors[251:250] = RED;
square ray_126(126,100 + ((MAX_HEIGHT - 167) / 2),1,167, x_pixel, y_pixel, is_in_rays[126]);
assign ray_colors[253:252] = RED;
square ray_127(127,100 + ((MAX_HEIGHT - 166) / 2),1,166, x_pixel, y_pixel, is_in_rays[127]);
assign ray_colors[255:254] = RED;
square ray_128(128,100 + ((MAX_HEIGHT - 165) / 2),1,165, x_pixel, y_pixel, is_in_rays[128]);
assign ray_colors[257:256] = RED;
square ray_129(129,100 + ((MAX_HEIGHT - 164) / 2),1,164, x_pixel, y_pixel, is_in_rays[129]);
assign ray_colors[259:258] = RED;
square ray_130(130,100 + ((MAX_HEIGHT - 164) / 2),1,164, x_pixel, y_pixel, is_in_rays[130]);
assign ray_colors[261:260] = RED;
square ray_131(131,100 + ((MAX_HEIGHT - 163) / 2),1,163, x_pixel, y_pixel, is_in_rays[131]);
assign ray_colors[263:262] = RED;
square ray_132(132,100 + ((MAX_HEIGHT - 162) / 2),1,162, x_pixel, y_pixel, is_in_rays[132]);
assign ray_colors[265:264] = RED;
square ray_133(133,100 + ((MAX_HEIGHT - 161) / 2),1,161, x_pixel, y_pixel, is_in_rays[133]);
assign ray_colors[267:266] = RED;
square ray_134(134,100 + ((MAX_HEIGHT - 160) / 2),1,160, x_pixel, y_pixel, is_in_rays[134]);
assign ray_colors[269:268] = RED;
square ray_135(135,100 + ((MAX_HEIGHT - 159) / 2),1,159, x_pixel, y_pixel, is_in_rays[135]);
assign ray_colors[271:270] = RED;
square ray_136(136,100 + ((MAX_HEIGHT - 159) / 2),1,159, x_pixel, y_pixel, is_in_rays[136]);
assign ray_colors[273:272] = RED;
square ray_137(137,100 + ((MAX_HEIGHT - 158) / 2),1,158, x_pixel, y_pixel, is_in_rays[137]);
assign ray_colors[275:274] = RED;
square ray_138(138,100 + ((MAX_HEIGHT - 157) / 2),1,157, x_pixel, y_pixel, is_in_rays[138]);
assign ray_colors[277:276] = RED;
square ray_139(139,100 + ((MAX_HEIGHT - 156) / 2),1,156, x_pixel, y_pixel, is_in_rays[139]);
assign ray_colors[279:278] = RED;
square ray_140(140,100 + ((MAX_HEIGHT - 155) / 2),1,155, x_pixel, y_pixel, is_in_rays[140]);
assign ray_colors[281:280] = RED;
square ray_141(141,100 + ((MAX_HEIGHT - 154) / 2),1,154, x_pixel, y_pixel, is_in_rays[141]);
assign ray_colors[283:282] = RED;
square ray_142(142,100 + ((MAX_HEIGHT - 153) / 2),1,153, x_pixel, y_pixel, is_in_rays[142]);
assign ray_colors[285:284] = RED;
square ray_143(143,100 + ((MAX_HEIGHT - 153) / 2),1,153, x_pixel, y_pixel, is_in_rays[143]);
assign ray_colors[287:286] = RED;
square ray_144(144,100 + ((MAX_HEIGHT - 152) / 2),1,152, x_pixel, y_pixel, is_in_rays[144]);
assign ray_colors[289:288] = RED;
square ray_145(145,100 + ((MAX_HEIGHT - 151) / 2),1,151, x_pixel, y_pixel, is_in_rays[145]);
assign ray_colors[291:290] = RED;
square ray_146(146,100 + ((MAX_HEIGHT - 150) / 2),1,150, x_pixel, y_pixel, is_in_rays[146]);
assign ray_colors[293:292] = RED;
square ray_147(147,100 + ((MAX_HEIGHT - 149) / 2),1,149, x_pixel, y_pixel, is_in_rays[147]);
assign ray_colors[295:294] = RED;
square ray_148(148,100 + ((MAX_HEIGHT - 148) / 2),1,148, x_pixel, y_pixel, is_in_rays[148]);
assign ray_colors[297:296] = RED;
square ray_149(149,100 + ((MAX_HEIGHT - 147) / 2),1,147, x_pixel, y_pixel, is_in_rays[149]);
assign ray_colors[299:298] = RED;
square ray_150(150,100 + ((MAX_HEIGHT - 147) / 2),1,147, x_pixel, y_pixel, is_in_rays[150]);
assign ray_colors[301:300] = RED;
square ray_151(151,100 + ((MAX_HEIGHT - 146) / 2),1,146, x_pixel, y_pixel, is_in_rays[151]);
assign ray_colors[303:302] = RED;
square ray_152(152,100 + ((MAX_HEIGHT - 145) / 2),1,145, x_pixel, y_pixel, is_in_rays[152]);
assign ray_colors[305:304] = RED;
square ray_153(153,100 + ((MAX_HEIGHT - 144) / 2),1,144, x_pixel, y_pixel, is_in_rays[153]);
assign ray_colors[307:306] = RED;
square ray_154(154,100 + ((MAX_HEIGHT - 143) / 2),1,143, x_pixel, y_pixel, is_in_rays[154]);
assign ray_colors[309:308] = RED;
square ray_155(155,100 + ((MAX_HEIGHT - 142) / 2),1,142, x_pixel, y_pixel, is_in_rays[155]);
assign ray_colors[311:310] = RED;
square ray_156(156,100 + ((MAX_HEIGHT - 141) / 2),1,141, x_pixel, y_pixel, is_in_rays[156]);
assign ray_colors[313:312] = RED;
square ray_157(157,100 + ((MAX_HEIGHT - 141) / 2),1,141, x_pixel, y_pixel, is_in_rays[157]);
assign ray_colors[315:314] = RED;
square ray_158(158,100 + ((MAX_HEIGHT - 140) / 2),1,140, x_pixel, y_pixel, is_in_rays[158]);
assign ray_colors[317:316] = RED;
square ray_159(159,100 + ((MAX_HEIGHT - 139) / 2),1,139, x_pixel, y_pixel, is_in_rays[159]);
assign ray_colors[319:318] = RED;
square ray_160(160,100 + ((MAX_HEIGHT - 138) / 2),1,138, x_pixel, y_pixel, is_in_rays[160]);
assign ray_colors[321:320] = RED;
square ray_161(161,100 + ((MAX_HEIGHT - 137) / 2),1,137, x_pixel, y_pixel, is_in_rays[161]);
assign ray_colors[323:322] = RED;
square ray_162(162,100 + ((MAX_HEIGHT - 136) / 2),1,136, x_pixel, y_pixel, is_in_rays[162]);
assign ray_colors[325:324] = RED;
square ray_163(163,100 + ((MAX_HEIGHT - 136) / 2),1,136, x_pixel, y_pixel, is_in_rays[163]);
assign ray_colors[327:326] = RED;
square ray_164(164,100 + ((MAX_HEIGHT - 135) / 2),1,135, x_pixel, y_pixel, is_in_rays[164]);
assign ray_colors[329:328] = RED;
square ray_165(165,100 + ((MAX_HEIGHT - 134) / 2),1,134, x_pixel, y_pixel, is_in_rays[165]);
assign ray_colors[331:330] = RED;
square ray_166(166,100 + ((MAX_HEIGHT - 133) / 2),1,133, x_pixel, y_pixel, is_in_rays[166]);
assign ray_colors[333:332] = RED;
square ray_167(167,100 + ((MAX_HEIGHT - 132) / 2),1,132, x_pixel, y_pixel, is_in_rays[167]);
assign ray_colors[335:334] = RED;
square ray_168(168,100 + ((MAX_HEIGHT - 131) / 2),1,131, x_pixel, y_pixel, is_in_rays[168]);
assign ray_colors[337:336] = RED;
square ray_169(169,100 + ((MAX_HEIGHT - 130) / 2),1,130, x_pixel, y_pixel, is_in_rays[169]);
assign ray_colors[339:338] = RED;
square ray_170(170,100 + ((MAX_HEIGHT - 130) / 2),1,130, x_pixel, y_pixel, is_in_rays[170]);
assign ray_colors[341:340] = RED;
square ray_171(171,100 + ((MAX_HEIGHT - 129) / 2),1,129, x_pixel, y_pixel, is_in_rays[171]);
assign ray_colors[343:342] = RED;
square ray_172(172,100 + ((MAX_HEIGHT - 128) / 2),1,128, x_pixel, y_pixel, is_in_rays[172]);
assign ray_colors[345:344] = RED;
square ray_173(173,100 + ((MAX_HEIGHT - 127) / 2),1,127, x_pixel, y_pixel, is_in_rays[173]);
assign ray_colors[347:346] = RED;
square ray_174(174,100 + ((MAX_HEIGHT - 126) / 2),1,126, x_pixel, y_pixel, is_in_rays[174]);
assign ray_colors[349:348] = RED;
square ray_175(175,100 + ((MAX_HEIGHT - 125) / 2),1,125, x_pixel, y_pixel, is_in_rays[175]);
assign ray_colors[351:350] = RED;
square ray_176(176,100 + ((MAX_HEIGHT - 124) / 2),1,124, x_pixel, y_pixel, is_in_rays[176]);
assign ray_colors[353:352] = RED;
square ray_177(177,100 + ((MAX_HEIGHT - 124) / 2),1,124, x_pixel, y_pixel, is_in_rays[177]);
assign ray_colors[355:354] = RED;
square ray_178(178,100 + ((MAX_HEIGHT - 123) / 2),1,123, x_pixel, y_pixel, is_in_rays[178]);
assign ray_colors[357:356] = RED;
square ray_179(179,100 + ((MAX_HEIGHT - 122) / 2),1,122, x_pixel, y_pixel, is_in_rays[179]);
assign ray_colors[359:358] = RED;
square ray_180(180,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[180]);
assign ray_colors[361:360] = BLUE;
square ray_181(181,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[181]);
assign ray_colors[363:362] = BLUE;
square ray_182(182,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[182]);
assign ray_colors[365:364] = BLUE;
square ray_183(183,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[183]);
assign ray_colors[367:366] = BLUE;
square ray_184(184,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[184]);
assign ray_colors[369:368] = BLUE;
square ray_185(185,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[185]);
assign ray_colors[371:370] = BLUE;
square ray_186(186,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[186]);
assign ray_colors[373:372] = BLUE;
square ray_187(187,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[187]);
assign ray_colors[375:374] = BLUE;
square ray_188(188,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[188]);
assign ray_colors[377:376] = BLUE;
square ray_189(189,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[189]);
assign ray_colors[379:378] = BLUE;
square ray_190(190,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[190]);
assign ray_colors[381:380] = BLUE;
square ray_191(191,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[191]);
assign ray_colors[383:382] = BLUE;
square ray_192(192,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[192]);
assign ray_colors[385:384] = BLUE;
square ray_193(193,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[193]);
assign ray_colors[387:386] = BLUE;
square ray_194(194,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[194]);
assign ray_colors[389:388] = BLUE;
square ray_195(195,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[195]);
assign ray_colors[391:390] = BLUE;
square ray_196(196,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[196]);
assign ray_colors[393:392] = BLUE;
square ray_197(197,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[197]);
assign ray_colors[395:394] = BLUE;
square ray_198(198,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[198]);
assign ray_colors[397:396] = BLUE;
square ray_199(199,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[199]);
assign ray_colors[399:398] = BLUE;
square ray_200(200,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[200]);
assign ray_colors[401:400] = BLUE;
square ray_201(201,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[201]);
assign ray_colors[403:402] = BLUE;
square ray_202(202,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[202]);
assign ray_colors[405:404] = BLUE;
square ray_203(203,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[203]);
assign ray_colors[407:406] = BLUE;
square ray_204(204,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[204]);
assign ray_colors[409:408] = BLUE;
square ray_205(205,100 + ((MAX_HEIGHT - 73) / 2),1,73, x_pixel, y_pixel, is_in_rays[205]);
assign ray_colors[411:410] = BLUE;
square ray_206(206,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[206]);
assign ray_colors[413:412] = BLUE;
square ray_207(207,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[207]);
assign ray_colors[415:414] = BLUE;
square ray_208(208,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[208]);
assign ray_colors[417:416] = BLUE;
square ray_209(209,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[209]);
assign ray_colors[419:418] = BLUE;
square ray_210(210,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[210]);
assign ray_colors[421:420] = BLUE;
square ray_211(211,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[211]);
assign ray_colors[423:422] = BLUE;
square ray_212(212,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[212]);
assign ray_colors[425:424] = BLUE;
square ray_213(213,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[213]);
assign ray_colors[427:426] = BLUE;
square ray_214(214,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[214]);
assign ray_colors[429:428] = BLUE;
square ray_215(215,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[215]);
assign ray_colors[431:430] = BLUE;
square ray_216(216,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[216]);
assign ray_colors[433:432] = BLUE;
square ray_217(217,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[217]);
assign ray_colors[435:434] = BLUE;
square ray_218(218,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[218]);
assign ray_colors[437:436] = BLUE;
square ray_219(219,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[219]);
assign ray_colors[439:438] = BLUE;
square ray_220(220,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[220]);
assign ray_colors[441:440] = BLUE;
square ray_221(221,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[221]);
assign ray_colors[443:442] = BLUE;
square ray_222(222,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[222]);
assign ray_colors[445:444] = BLUE;
square ray_223(223,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[223]);
assign ray_colors[447:446] = BLUE;
square ray_224(224,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[224]);
assign ray_colors[449:448] = BLUE;
square ray_225(225,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[225]);
assign ray_colors[451:450] = BLUE;
square ray_226(226,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[226]);
assign ray_colors[453:452] = BLUE;
square ray_227(227,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[227]);
assign ray_colors[455:454] = BLUE;
square ray_228(228,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[228]);
assign ray_colors[457:456] = BLUE;
square ray_229(229,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[229]);
assign ray_colors[459:458] = BLUE;
square ray_230(230,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[230]);
assign ray_colors[461:460] = BLUE;
square ray_231(231,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[231]);
assign ray_colors[463:462] = BLUE;
square ray_232(232,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[232]);
assign ray_colors[465:464] = BLUE;
square ray_233(233,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[233]);
assign ray_colors[467:466] = BLUE;
square ray_234(234,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[234]);
assign ray_colors[469:468] = BLUE;
square ray_235(235,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[235]);
assign ray_colors[471:470] = BLUE;
square ray_236(236,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[236]);
assign ray_colors[473:472] = BLUE;
square ray_237(237,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[237]);
assign ray_colors[475:474] = BLUE;
square ray_238(238,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[238]);
assign ray_colors[477:476] = BLUE;
square ray_239(239,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[239]);
assign ray_colors[479:478] = BLUE;
square ray_240(240,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[240]);
assign ray_colors[481:480] = BLUE;
square ray_241(241,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[241]);
assign ray_colors[483:482] = BLUE;
square ray_242(242,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[242]);
assign ray_colors[485:484] = BLUE;
square ray_243(243,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[243]);
assign ray_colors[487:486] = BLUE;
square ray_244(244,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[244]);
assign ray_colors[489:488] = BLUE;
square ray_245(245,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[245]);
assign ray_colors[491:490] = BLUE;
square ray_246(246,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[246]);
assign ray_colors[493:492] = BLUE;
square ray_247(247,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[247]);
assign ray_colors[495:494] = BLUE;
square ray_248(248,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[248]);
assign ray_colors[497:496] = BLUE;
square ray_249(249,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[249]);
assign ray_colors[499:498] = BLUE;
square ray_250(250,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[250]);
assign ray_colors[501:500] = BLUE;
square ray_251(251,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[251]);
assign ray_colors[503:502] = BLUE;
square ray_252(252,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[252]);
assign ray_colors[505:504] = BLUE;
square ray_253(253,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[253]);
assign ray_colors[507:506] = BLUE;
square ray_254(254,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[254]);
assign ray_colors[509:508] = BLUE;
square ray_255(255,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[255]);
assign ray_colors[511:510] = BLUE;
square ray_256(256,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[256]);
assign ray_colors[513:512] = BLUE;
square ray_257(257,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[257]);
assign ray_colors[515:514] = BLUE;
square ray_258(258,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[258]);
assign ray_colors[517:516] = BLUE;
square ray_259(259,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[259]);
assign ray_colors[519:518] = BLUE;
square ray_260(260,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[260]);
assign ray_colors[521:520] = BLUE;
square ray_261(261,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[261]);
assign ray_colors[523:522] = BLUE;
square ray_262(262,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[262]);
assign ray_colors[525:524] = BLUE;
square ray_263(263,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[263]);
assign ray_colors[527:526] = BLUE;
square ray_264(264,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[264]);
assign ray_colors[529:528] = BLUE;
square ray_265(265,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[265]);
assign ray_colors[531:530] = BLUE;
square ray_266(266,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[266]);
assign ray_colors[533:532] = BLUE;
square ray_267(267,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[267]);
assign ray_colors[535:534] = BLUE;
square ray_268(268,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[268]);
assign ray_colors[537:536] = BLUE;
square ray_269(269,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[269]);
assign ray_colors[539:538] = BLUE;
square ray_270(270,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[270]);
assign ray_colors[541:540] = BLUE;
square ray_271(271,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[271]);
assign ray_colors[543:542] = BLUE;
square ray_272(272,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[272]);
assign ray_colors[545:544] = BLUE;
square ray_273(273,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[273]);
assign ray_colors[547:546] = BLUE;
square ray_274(274,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[274]);
assign ray_colors[549:548] = BLUE;
square ray_275(275,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[275]);
assign ray_colors[551:550] = BLUE;
square ray_276(276,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[276]);
assign ray_colors[553:552] = BLUE;
square ray_277(277,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[277]);
assign ray_colors[555:554] = BLUE;
square ray_278(278,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[278]);
assign ray_colors[557:556] = BLUE;
square ray_279(279,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[279]);
assign ray_colors[559:558] = BLUE;
square ray_280(280,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[280]);
assign ray_colors[561:560] = BLUE;
square ray_281(281,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[281]);
assign ray_colors[563:562] = BLUE;
square ray_282(282,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[282]);
assign ray_colors[565:564] = BLUE;
square ray_283(283,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[283]);
assign ray_colors[567:566] = BLUE;
square ray_284(284,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[284]);
assign ray_colors[569:568] = BLUE;
square ray_285(285,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[285]);
assign ray_colors[571:570] = BLUE;
square ray_286(286,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[286]);
assign ray_colors[573:572] = BLUE;
square ray_287(287,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[287]);
assign ray_colors[575:574] = BLUE;
square ray_288(288,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[288]);
assign ray_colors[577:576] = BLUE;
square ray_289(289,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[289]);
assign ray_colors[579:578] = BLUE;
square ray_290(290,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[290]);
assign ray_colors[581:580] = BLUE;
square ray_291(291,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[291]);
assign ray_colors[583:582] = BLUE;
square ray_292(292,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[292]);
assign ray_colors[585:584] = BLUE;
square ray_293(293,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[293]);
assign ray_colors[587:586] = BLUE;
square ray_294(294,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[294]);
assign ray_colors[589:588] = BLUE;
square ray_295(295,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[295]);
assign ray_colors[591:590] = BLUE;
square ray_296(296,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[296]);
assign ray_colors[593:592] = BLUE;
square ray_297(297,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[297]);
assign ray_colors[595:594] = BLUE;
square ray_298(298,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[298]);
assign ray_colors[597:596] = BLUE;
square ray_299(299,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[299]);
assign ray_colors[599:598] = BLUE;
square ray_300(300,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[300]);
assign ray_colors[601:600] = BLUE;
square ray_301(301,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[301]);
assign ray_colors[603:602] = BLUE;
square ray_302(302,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[302]);
assign ray_colors[605:604] = BLUE;
square ray_303(303,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[303]);
assign ray_colors[607:606] = BLUE;
square ray_304(304,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[304]);
assign ray_colors[609:608] = BLUE;
square ray_305(305,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[305]);
assign ray_colors[611:610] = BLUE;
square ray_306(306,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[306]);
assign ray_colors[613:612] = BLUE;
square ray_307(307,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[307]);
assign ray_colors[615:614] = BLUE;
square ray_308(308,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[308]);
assign ray_colors[617:616] = BLUE;
square ray_309(309,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[309]);
assign ray_colors[619:618] = BLUE;
square ray_310(310,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[310]);
assign ray_colors[621:620] = BLUE;
square ray_311(311,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[311]);
assign ray_colors[623:622] = BLUE;
square ray_312(312,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[312]);
assign ray_colors[625:624] = BLUE;
square ray_313(313,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[313]);
assign ray_colors[627:626] = BLUE;
square ray_314(314,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[314]);
assign ray_colors[629:628] = BLUE;
square ray_315(315,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[315]);
assign ray_colors[631:630] = BLUE;
square ray_316(316,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[316]);
assign ray_colors[633:632] = BLUE;
square ray_317(317,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[317]);
assign ray_colors[635:634] = BLUE;
square ray_318(318,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[318]);
assign ray_colors[637:636] = BLUE;
square ray_319(319,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[319]);
assign ray_colors[639:638] = BLUE;
square ray_320(320,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[320]);
assign ray_colors[641:640] = BLUE;
square ray_321(321,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[321]);
assign ray_colors[643:642] = BLUE;
square ray_322(322,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[322]);
assign ray_colors[645:644] = BLUE;
square ray_323(323,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[323]);
assign ray_colors[647:646] = BLUE;
square ray_324(324,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[324]);
assign ray_colors[649:648] = BLUE;
square ray_325(325,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[325]);
assign ray_colors[651:650] = BLUE;
square ray_326(326,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[326]);
assign ray_colors[653:652] = BLUE;
square ray_327(327,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[327]);
assign ray_colors[655:654] = BLUE;
square ray_328(328,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[328]);
assign ray_colors[657:656] = BLUE;
square ray_329(329,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[329]);
assign ray_colors[659:658] = BLUE;
square ray_330(330,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[330]);
assign ray_colors[661:660] = BLUE;
square ray_331(331,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[331]);
assign ray_colors[663:662] = BLUE;
square ray_332(332,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[332]);
assign ray_colors[665:664] = BLUE;
square ray_333(333,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[333]);
assign ray_colors[667:666] = BLUE;
square ray_334(334,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[334]);
assign ray_colors[669:668] = BLUE;
square ray_335(335,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[335]);
assign ray_colors[671:670] = BLUE;
square ray_336(336,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[336]);
assign ray_colors[673:672] = BLUE;
square ray_337(337,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[337]);
assign ray_colors[675:674] = BLUE;
square ray_338(338,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[338]);
assign ray_colors[677:676] = BLUE;
square ray_339(339,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[339]);
assign ray_colors[679:678] = BLUE;
square ray_340(340,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[340]);
assign ray_colors[681:680] = BLUE;
square ray_341(341,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[341]);
assign ray_colors[683:682] = BLUE;
square ray_342(342,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[342]);
assign ray_colors[685:684] = BLUE;
square ray_343(343,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[343]);
assign ray_colors[687:686] = BLUE;
square ray_344(344,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[344]);
assign ray_colors[689:688] = BLUE;
square ray_345(345,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[345]);
assign ray_colors[691:690] = BLUE;
square ray_346(346,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[346]);
assign ray_colors[693:692] = BLUE;
square ray_347(347,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[347]);
assign ray_colors[695:694] = BLUE;
square ray_348(348,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[348]);
assign ray_colors[697:696] = BLUE;
square ray_349(349,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[349]);
assign ray_colors[699:698] = BLUE;
square ray_350(350,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[350]);
assign ray_colors[701:700] = BLUE;
square ray_351(351,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[351]);
assign ray_colors[703:702] = BLUE;
square ray_352(352,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[352]);
assign ray_colors[705:704] = BLUE;
square ray_353(353,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[353]);
assign ray_colors[707:706] = BLUE;
square ray_354(354,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[354]);
assign ray_colors[709:708] = BLUE;
square ray_355(355,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[355]);
assign ray_colors[711:710] = BLUE;
square ray_356(356,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[356]);
assign ray_colors[713:712] = BLUE;
square ray_357(357,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[357]);
assign ray_colors[715:714] = BLUE;
square ray_358(358,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[358]);
assign ray_colors[717:716] = BLUE;
square ray_359(359,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[359]);
assign ray_colors[719:718] = BLUE;
square ray_360(360,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[360]);
assign ray_colors[721:720] = BLUE;
square ray_361(361,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[361]);
assign ray_colors[723:722] = BLUE;
square ray_362(362,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[362]);
assign ray_colors[725:724] = BLUE;
square ray_363(363,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[363]);
assign ray_colors[727:726] = BLUE;
square ray_364(364,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[364]);
assign ray_colors[729:728] = BLUE;
square ray_365(365,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[365]);
assign ray_colors[731:730] = BLUE;
square ray_366(366,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[366]);
assign ray_colors[733:732] = BLUE;
square ray_367(367,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[367]);
assign ray_colors[735:734] = BLUE;
square ray_368(368,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[368]);
assign ray_colors[737:736] = BLUE;
square ray_369(369,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[369]);
assign ray_colors[739:738] = BLUE;
square ray_370(370,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[370]);
assign ray_colors[741:740] = BLUE;
square ray_371(371,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[371]);
assign ray_colors[743:742] = BLUE;
square ray_372(372,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[372]);
assign ray_colors[745:744] = BLUE;
square ray_373(373,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[373]);
assign ray_colors[747:746] = BLUE;
square ray_374(374,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[374]);
assign ray_colors[749:748] = BLUE;
square ray_375(375,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[375]);
assign ray_colors[751:750] = BLUE;
square ray_376(376,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[376]);
assign ray_colors[753:752] = BLUE;
square ray_377(377,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[377]);
assign ray_colors[755:754] = BLUE;
square ray_378(378,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[378]);
assign ray_colors[757:756] = BLUE;
square ray_379(379,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[379]);
assign ray_colors[759:758] = BLUE;
square ray_380(380,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[380]);
assign ray_colors[761:760] = BLUE;
square ray_381(381,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[381]);
assign ray_colors[763:762] = BLUE;
square ray_382(382,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[382]);
assign ray_colors[765:764] = BLUE;
square ray_383(383,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[383]);
assign ray_colors[767:766] = BLUE;
square ray_384(384,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[384]);
assign ray_colors[769:768] = BLUE;
square ray_385(385,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[385]);
assign ray_colors[771:770] = BLUE;
square ray_386(386,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[386]);
assign ray_colors[773:772] = BLUE;
square ray_387(387,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[387]);
assign ray_colors[775:774] = BLUE;
square ray_388(388,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[388]);
assign ray_colors[777:776] = BLUE;
square ray_389(389,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[389]);
assign ray_colors[779:778] = BLUE;
square ray_390(390,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[390]);
assign ray_colors[781:780] = BLUE;
square ray_391(391,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[391]);
assign ray_colors[783:782] = BLUE;
square ray_392(392,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[392]);
assign ray_colors[785:784] = BLUE;
square ray_393(393,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[393]);
assign ray_colors[787:786] = BLUE;
square ray_394(394,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[394]);
assign ray_colors[789:788] = BLUE;
square ray_395(395,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[395]);
assign ray_colors[791:790] = BLUE;
square ray_396(396,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[396]);
assign ray_colors[793:792] = BLUE;
square ray_397(397,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[397]);
assign ray_colors[795:794] = BLUE;
square ray_398(398,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[398]);
assign ray_colors[797:796] = BLUE;
square ray_399(399,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[399]);
assign ray_colors[799:798] = BLUE;
square ray_400(400,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[400]);
assign ray_colors[801:800] = BLUE;
square ray_401(401,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[401]);
assign ray_colors[803:802] = BLUE;
square ray_402(402,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[402]);
assign ray_colors[805:804] = BLUE;
square ray_403(403,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[403]);
assign ray_colors[807:806] = BLUE;
square ray_404(404,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[404]);
assign ray_colors[809:808] = BLUE;
square ray_405(405,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[405]);
assign ray_colors[811:810] = BLUE;
square ray_406(406,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[406]);
assign ray_colors[813:812] = BLUE;
square ray_407(407,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[407]);
assign ray_colors[815:814] = BLUE;
square ray_408(408,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[408]);
assign ray_colors[817:816] = BLUE;
square ray_409(409,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[409]);
assign ray_colors[819:818] = BLUE;
square ray_410(410,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[410]);
assign ray_colors[821:820] = BLUE;
square ray_411(411,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[411]);
assign ray_colors[823:822] = BLUE;
square ray_412(412,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[412]);
assign ray_colors[825:824] = BLUE;
square ray_413(413,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[413]);
assign ray_colors[827:826] = BLUE;
square ray_414(414,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[414]);
assign ray_colors[829:828] = BLUE;
square ray_415(415,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[415]);
assign ray_colors[831:830] = BLUE;
square ray_416(416,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[416]);
assign ray_colors[833:832] = BLUE;
square ray_417(417,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[417]);
assign ray_colors[835:834] = BLUE;
square ray_418(418,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[418]);
assign ray_colors[837:836] = BLUE;
square ray_419(419,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[419]);
assign ray_colors[839:838] = BLUE;
square ray_420(420,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[420]);
assign ray_colors[841:840] = BLUE;
square ray_421(421,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[421]);
assign ray_colors[843:842] = BLUE;
square ray_422(422,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[422]);
assign ray_colors[845:844] = BLUE;
square ray_423(423,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[423]);
assign ray_colors[847:846] = BLUE;
square ray_424(424,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[424]);
assign ray_colors[849:848] = BLUE;
square ray_425(425,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[425]);
assign ray_colors[851:850] = BLUE;
square ray_426(426,100 + ((MAX_HEIGHT - 74) / 2),1,74, x_pixel, y_pixel, is_in_rays[426]);
assign ray_colors[853:852] = BLUE;
square ray_427(427,100 + ((MAX_HEIGHT - 93) / 2),1,93, x_pixel, y_pixel, is_in_rays[427]);
assign ray_colors[855:854] = GREEN;
square ray_428(428,100 + ((MAX_HEIGHT - 93) / 2),1,93, x_pixel, y_pixel, is_in_rays[428]);
assign ray_colors[857:856] = GREEN;
square ray_429(429,100 + ((MAX_HEIGHT - 94) / 2),1,94, x_pixel, y_pixel, is_in_rays[429]);
assign ray_colors[859:858] = GREEN;
square ray_430(430,100 + ((MAX_HEIGHT - 95) / 2),1,95, x_pixel, y_pixel, is_in_rays[430]);
assign ray_colors[861:860] = GREEN;
square ray_431(431,100 + ((MAX_HEIGHT - 96) / 2),1,96, x_pixel, y_pixel, is_in_rays[431]);
assign ray_colors[863:862] = GREEN;
square ray_432(432,100 + ((MAX_HEIGHT - 97) / 2),1,97, x_pixel, y_pixel, is_in_rays[432]);
assign ray_colors[865:864] = GREEN;
square ray_433(433,100 + ((MAX_HEIGHT - 98) / 2),1,98, x_pixel, y_pixel, is_in_rays[433]);
assign ray_colors[867:866] = GREEN;
square ray_434(434,100 + ((MAX_HEIGHT - 99) / 2),1,99, x_pixel, y_pixel, is_in_rays[434]);
assign ray_colors[869:868] = GREEN;
square ray_435(435,100 + ((MAX_HEIGHT - 99) / 2),1,99, x_pixel, y_pixel, is_in_rays[435]);
assign ray_colors[871:870] = GREEN;
square ray_436(436,100 + ((MAX_HEIGHT - 100) / 2),1,100, x_pixel, y_pixel, is_in_rays[436]);
assign ray_colors[873:872] = GREEN;
square ray_437(437,100 + ((MAX_HEIGHT - 101) / 2),1,101, x_pixel, y_pixel, is_in_rays[437]);
assign ray_colors[875:874] = GREEN;
square ray_438(438,100 + ((MAX_HEIGHT - 102) / 2),1,102, x_pixel, y_pixel, is_in_rays[438]);
assign ray_colors[877:876] = GREEN;
square ray_439(439,100 + ((MAX_HEIGHT - 103) / 2),1,103, x_pixel, y_pixel, is_in_rays[439]);
assign ray_colors[879:878] = GREEN;
square ray_440(440,100 + ((MAX_HEIGHT - 104) / 2),1,104, x_pixel, y_pixel, is_in_rays[440]);
assign ray_colors[881:880] = GREEN;
square ray_441(441,100 + ((MAX_HEIGHT - 105) / 2),1,105, x_pixel, y_pixel, is_in_rays[441]);
assign ray_colors[883:882] = GREEN;
square ray_442(442,100 + ((MAX_HEIGHT - 106) / 2),1,106, x_pixel, y_pixel, is_in_rays[442]);
assign ray_colors[885:884] = GREEN;
square ray_443(443,100 + ((MAX_HEIGHT - 106) / 2),1,106, x_pixel, y_pixel, is_in_rays[443]);
assign ray_colors[887:886] = GREEN;
square ray_444(444,100 + ((MAX_HEIGHT - 107) / 2),1,107, x_pixel, y_pixel, is_in_rays[444]);
assign ray_colors[889:888] = GREEN;
square ray_445(445,100 + ((MAX_HEIGHT - 108) / 2),1,108, x_pixel, y_pixel, is_in_rays[445]);
assign ray_colors[891:890] = GREEN;
square ray_446(446,100 + ((MAX_HEIGHT - 109) / 2),1,109, x_pixel, y_pixel, is_in_rays[446]);
assign ray_colors[893:892] = GREEN;
square ray_447(447,100 + ((MAX_HEIGHT - 110) / 2),1,110, x_pixel, y_pixel, is_in_rays[447]);
assign ray_colors[895:894] = GREEN;
square ray_448(448,100 + ((MAX_HEIGHT - 111) / 2),1,111, x_pixel, y_pixel, is_in_rays[448]);
assign ray_colors[897:896] = GREEN;
square ray_449(449,100 + ((MAX_HEIGHT - 112) / 2),1,112, x_pixel, y_pixel, is_in_rays[449]);
assign ray_colors[899:898] = GREEN;
square ray_450(450,100 + ((MAX_HEIGHT - 112) / 2),1,112, x_pixel, y_pixel, is_in_rays[450]);
assign ray_colors[901:900] = GREEN;
square ray_451(451,100 + ((MAX_HEIGHT - 113) / 2),1,113, x_pixel, y_pixel, is_in_rays[451]);
assign ray_colors[903:902] = GREEN;
square ray_452(452,100 + ((MAX_HEIGHT - 114) / 2),1,114, x_pixel, y_pixel, is_in_rays[452]);
assign ray_colors[905:904] = GREEN;
square ray_453(453,100 + ((MAX_HEIGHT - 115) / 2),1,115, x_pixel, y_pixel, is_in_rays[453]);
assign ray_colors[907:906] = GREEN;
square ray_454(454,100 + ((MAX_HEIGHT - 116) / 2),1,116, x_pixel, y_pixel, is_in_rays[454]);
assign ray_colors[909:908] = GREEN;
square ray_455(455,100 + ((MAX_HEIGHT - 117) / 2),1,117, x_pixel, y_pixel, is_in_rays[455]);
assign ray_colors[911:910] = GREEN;
square ray_456(456,100 + ((MAX_HEIGHT - 118) / 2),1,118, x_pixel, y_pixel, is_in_rays[456]);
assign ray_colors[913:912] = GREEN;
square ray_457(457,100 + ((MAX_HEIGHT - 118) / 2),1,118, x_pixel, y_pixel, is_in_rays[457]);
assign ray_colors[915:914] = GREEN;
square ray_458(458,100 + ((MAX_HEIGHT - 119) / 2),1,119, x_pixel, y_pixel, is_in_rays[458]);
assign ray_colors[917:916] = GREEN;
square ray_459(459,100 + ((MAX_HEIGHT - 120) / 2),1,120, x_pixel, y_pixel, is_in_rays[459]);
assign ray_colors[919:918] = GREEN;
square ray_460(460,100 + ((MAX_HEIGHT - 121) / 2),1,121, x_pixel, y_pixel, is_in_rays[460]);
assign ray_colors[921:920] = GREEN;
square ray_461(461,100 + ((MAX_HEIGHT - 122) / 2),1,122, x_pixel, y_pixel, is_in_rays[461]);
assign ray_colors[923:922] = GREEN;
square ray_462(462,100 + ((MAX_HEIGHT - 123) / 2),1,123, x_pixel, y_pixel, is_in_rays[462]);
assign ray_colors[925:924] = GREEN;
square ray_463(463,100 + ((MAX_HEIGHT - 124) / 2),1,124, x_pixel, y_pixel, is_in_rays[463]);
assign ray_colors[927:926] = GREEN;
square ray_464(464,100 + ((MAX_HEIGHT - 124) / 2),1,124, x_pixel, y_pixel, is_in_rays[464]);
assign ray_colors[929:928] = GREEN;
square ray_465(465,100 + ((MAX_HEIGHT - 125) / 2),1,125, x_pixel, y_pixel, is_in_rays[465]);
assign ray_colors[931:930] = GREEN;
square ray_466(466,100 + ((MAX_HEIGHT - 126) / 2),1,126, x_pixel, y_pixel, is_in_rays[466]);
assign ray_colors[933:932] = GREEN;
square ray_467(467,100 + ((MAX_HEIGHT - 127) / 2),1,127, x_pixel, y_pixel, is_in_rays[467]);
assign ray_colors[935:934] = GREEN;
square ray_468(468,100 + ((MAX_HEIGHT - 128) / 2),1,128, x_pixel, y_pixel, is_in_rays[468]);
assign ray_colors[937:936] = GREEN;
square ray_469(469,100 + ((MAX_HEIGHT - 129) / 2),1,129, x_pixel, y_pixel, is_in_rays[469]);
assign ray_colors[939:938] = GREEN;
square ray_470(470,100 + ((MAX_HEIGHT - 130) / 2),1,130, x_pixel, y_pixel, is_in_rays[470]);
assign ray_colors[941:940] = GREEN;
square ray_471(471,100 + ((MAX_HEIGHT - 130) / 2),1,130, x_pixel, y_pixel, is_in_rays[471]);
assign ray_colors[943:942] = GREEN;
square ray_472(472,100 + ((MAX_HEIGHT - 131) / 2),1,131, x_pixel, y_pixel, is_in_rays[472]);
assign ray_colors[945:944] = GREEN;
square ray_473(473,100 + ((MAX_HEIGHT - 132) / 2),1,132, x_pixel, y_pixel, is_in_rays[473]);
assign ray_colors[947:946] = GREEN;
square ray_474(474,100 + ((MAX_HEIGHT - 133) / 2),1,133, x_pixel, y_pixel, is_in_rays[474]);
assign ray_colors[949:948] = GREEN;
square ray_475(475,100 + ((MAX_HEIGHT - 134) / 2),1,134, x_pixel, y_pixel, is_in_rays[475]);
assign ray_colors[951:950] = GREEN;
square ray_476(476,100 + ((MAX_HEIGHT - 135) / 2),1,135, x_pixel, y_pixel, is_in_rays[476]);
assign ray_colors[953:952] = GREEN;
square ray_477(477,100 + ((MAX_HEIGHT - 136) / 2),1,136, x_pixel, y_pixel, is_in_rays[477]);
assign ray_colors[955:954] = GREEN;
square ray_478(478,100 + ((MAX_HEIGHT - 136) / 2),1,136, x_pixel, y_pixel, is_in_rays[478]);
assign ray_colors[957:956] = GREEN;
square ray_479(479,100 + ((MAX_HEIGHT - 137) / 2),1,137, x_pixel, y_pixel, is_in_rays[479]);
assign ray_colors[959:958] = GREEN;
square ray_480(480,100 + ((MAX_HEIGHT - 138) / 2),1,138, x_pixel, y_pixel, is_in_rays[480]);
assign ray_colors[961:960] = GREEN;
square ray_481(481,100 + ((MAX_HEIGHT - 139) / 2),1,139, x_pixel, y_pixel, is_in_rays[481]);
assign ray_colors[963:962] = GREEN;
square ray_482(482,100 + ((MAX_HEIGHT - 140) / 2),1,140, x_pixel, y_pixel, is_in_rays[482]);
assign ray_colors[965:964] = GREEN;
square ray_483(483,100 + ((MAX_HEIGHT - 141) / 2),1,141, x_pixel, y_pixel, is_in_rays[483]);
assign ray_colors[967:966] = GREEN;
square ray_484(484,100 + ((MAX_HEIGHT - 141) / 2),1,141, x_pixel, y_pixel, is_in_rays[484]);
assign ray_colors[969:968] = GREEN;
square ray_485(485,100 + ((MAX_HEIGHT - 142) / 2),1,142, x_pixel, y_pixel, is_in_rays[485]);
assign ray_colors[971:970] = GREEN;
square ray_486(486,100 + ((MAX_HEIGHT - 143) / 2),1,143, x_pixel, y_pixel, is_in_rays[486]);
assign ray_colors[973:972] = GREEN;
square ray_487(487,100 + ((MAX_HEIGHT - 144) / 2),1,144, x_pixel, y_pixel, is_in_rays[487]);
assign ray_colors[975:974] = GREEN;
square ray_488(488,100 + ((MAX_HEIGHT - 145) / 2),1,145, x_pixel, y_pixel, is_in_rays[488]);
assign ray_colors[977:976] = GREEN;
square ray_489(489,100 + ((MAX_HEIGHT - 146) / 2),1,146, x_pixel, y_pixel, is_in_rays[489]);
assign ray_colors[979:978] = GREEN;
square ray_490(490,100 + ((MAX_HEIGHT - 147) / 2),1,147, x_pixel, y_pixel, is_in_rays[490]);
assign ray_colors[981:980] = GREEN;
square ray_491(491,100 + ((MAX_HEIGHT - 147) / 2),1,147, x_pixel, y_pixel, is_in_rays[491]);
assign ray_colors[983:982] = GREEN;
square ray_492(492,100 + ((MAX_HEIGHT - 148) / 2),1,148, x_pixel, y_pixel, is_in_rays[492]);
assign ray_colors[985:984] = GREEN;
square ray_493(493,100 + ((MAX_HEIGHT - 149) / 2),1,149, x_pixel, y_pixel, is_in_rays[493]);
assign ray_colors[987:986] = GREEN;
square ray_494(494,100 + ((MAX_HEIGHT - 150) / 2),1,150, x_pixel, y_pixel, is_in_rays[494]);
assign ray_colors[989:988] = GREEN;
square ray_495(495,100 + ((MAX_HEIGHT - 151) / 2),1,151, x_pixel, y_pixel, is_in_rays[495]);
assign ray_colors[991:990] = GREEN;
square ray_496(496,100 + ((MAX_HEIGHT - 152) / 2),1,152, x_pixel, y_pixel, is_in_rays[496]);
assign ray_colors[993:992] = GREEN;
square ray_497(497,100 + ((MAX_HEIGHT - 153) / 2),1,153, x_pixel, y_pixel, is_in_rays[497]);
assign ray_colors[995:994] = GREEN;
square ray_498(498,100 + ((MAX_HEIGHT - 153) / 2),1,153, x_pixel, y_pixel, is_in_rays[498]);
assign ray_colors[997:996] = GREEN;
square ray_499(499,100 + ((MAX_HEIGHT - 154) / 2),1,154, x_pixel, y_pixel, is_in_rays[499]);
assign ray_colors[999:998] = GREEN;
square ray_500(500,100 + ((MAX_HEIGHT - 155) / 2),1,155, x_pixel, y_pixel, is_in_rays[500]);
assign ray_colors[1001:1000] = GREEN;
square ray_501(501,100 + ((MAX_HEIGHT - 156) / 2),1,156, x_pixel, y_pixel, is_in_rays[501]);
assign ray_colors[1003:1002] = GREEN;
square ray_502(502,100 + ((MAX_HEIGHT - 157) / 2),1,157, x_pixel, y_pixel, is_in_rays[502]);
assign ray_colors[1005:1004] = GREEN;
square ray_503(503,100 + ((MAX_HEIGHT - 158) / 2),1,158, x_pixel, y_pixel, is_in_rays[503]);
assign ray_colors[1007:1006] = GREEN;
square ray_504(504,100 + ((MAX_HEIGHT - 159) / 2),1,159, x_pixel, y_pixel, is_in_rays[504]);
assign ray_colors[1009:1008] = GREEN;
square ray_505(505,100 + ((MAX_HEIGHT - 159) / 2),1,159, x_pixel, y_pixel, is_in_rays[505]);
assign ray_colors[1011:1010] = GREEN;
square ray_506(506,100 + ((MAX_HEIGHT - 160) / 2),1,160, x_pixel, y_pixel, is_in_rays[506]);
assign ray_colors[1013:1012] = GREEN;
square ray_507(507,100 + ((MAX_HEIGHT - 161) / 2),1,161, x_pixel, y_pixel, is_in_rays[507]);
assign ray_colors[1015:1014] = GREEN;
square ray_508(508,100 + ((MAX_HEIGHT - 162) / 2),1,162, x_pixel, y_pixel, is_in_rays[508]);
assign ray_colors[1017:1016] = GREEN;
square ray_509(509,100 + ((MAX_HEIGHT - 163) / 2),1,163, x_pixel, y_pixel, is_in_rays[509]);
assign ray_colors[1019:1018] = GREEN;
square ray_510(510,100 + ((MAX_HEIGHT - 164) / 2),1,164, x_pixel, y_pixel, is_in_rays[510]);
assign ray_colors[1021:1020] = GREEN;
square ray_511(511,100 + ((MAX_HEIGHT - 164) / 2),1,164, x_pixel, y_pixel, is_in_rays[511]);
assign ray_colors[1023:1022] = GREEN;
square ray_512(512,100 + ((MAX_HEIGHT - 165) / 2),1,165, x_pixel, y_pixel, is_in_rays[512]);
assign ray_colors[1025:1024] = GREEN;
square ray_513(513,100 + ((MAX_HEIGHT - 166) / 2),1,166, x_pixel, y_pixel, is_in_rays[513]);
assign ray_colors[1027:1026] = GREEN;
square ray_514(514,100 + ((MAX_HEIGHT - 167) / 2),1,167, x_pixel, y_pixel, is_in_rays[514]);
assign ray_colors[1029:1028] = GREEN;
square ray_515(515,100 + ((MAX_HEIGHT - 168) / 2),1,168, x_pixel, y_pixel, is_in_rays[515]);
assign ray_colors[1031:1030] = GREEN;
square ray_516(516,100 + ((MAX_HEIGHT - 169) / 2),1,169, x_pixel, y_pixel, is_in_rays[516]);
assign ray_colors[1033:1032] = GREEN;
square ray_517(517,100 + ((MAX_HEIGHT - 170) / 2),1,170, x_pixel, y_pixel, is_in_rays[517]);
assign ray_colors[1035:1034] = GREEN;
square ray_518(518,100 + ((MAX_HEIGHT - 170) / 2),1,170, x_pixel, y_pixel, is_in_rays[518]);
assign ray_colors[1037:1036] = GREEN;
square ray_519(519,100 + ((MAX_HEIGHT - 171) / 2),1,171, x_pixel, y_pixel, is_in_rays[519]);
assign ray_colors[1039:1038] = GREEN;
square ray_520(520,100 + ((MAX_HEIGHT - 172) / 2),1,172, x_pixel, y_pixel, is_in_rays[520]);
assign ray_colors[1041:1040] = GREEN;
square ray_521(521,100 + ((MAX_HEIGHT - 173) / 2),1,173, x_pixel, y_pixel, is_in_rays[521]);
assign ray_colors[1043:1042] = GREEN;
square ray_522(522,100 + ((MAX_HEIGHT - 174) / 2),1,174, x_pixel, y_pixel, is_in_rays[522]);
assign ray_colors[1045:1044] = GREEN;
square ray_523(523,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[523]);
assign ray_colors[1047:1046] = GREEN;
square ray_524(524,100 + ((MAX_HEIGHT - 175) / 2),1,175, x_pixel, y_pixel, is_in_rays[524]);
assign ray_colors[1049:1048] = GREEN;
square ray_525(525,100 + ((MAX_HEIGHT - 176) / 2),1,176, x_pixel, y_pixel, is_in_rays[525]);
assign ray_colors[1051:1050] = GREEN;
square ray_526(526,100 + ((MAX_HEIGHT - 177) / 2),1,177, x_pixel, y_pixel, is_in_rays[526]);
assign ray_colors[1053:1052] = GREEN;
square ray_527(527,100 + ((MAX_HEIGHT - 178) / 2),1,178, x_pixel, y_pixel, is_in_rays[527]);
assign ray_colors[1055:1054] = GREEN;
square ray_528(528,100 + ((MAX_HEIGHT - 179) / 2),1,179, x_pixel, y_pixel, is_in_rays[528]);
assign ray_colors[1057:1056] = GREEN;
square ray_529(529,100 + ((MAX_HEIGHT - 180) / 2),1,180, x_pixel, y_pixel, is_in_rays[529]);
assign ray_colors[1059:1058] = GREEN;
square ray_530(530,100 + ((MAX_HEIGHT - 181) / 2),1,181, x_pixel, y_pixel, is_in_rays[530]);
assign ray_colors[1061:1060] = GREEN;
square ray_531(531,100 + ((MAX_HEIGHT - 181) / 2),1,181, x_pixel, y_pixel, is_in_rays[531]);
assign ray_colors[1063:1062] = GREEN;
square ray_532(532,100 + ((MAX_HEIGHT - 182) / 2),1,182, x_pixel, y_pixel, is_in_rays[532]);
assign ray_colors[1065:1064] = GREEN;
square ray_533(533,100 + ((MAX_HEIGHT - 183) / 2),1,183, x_pixel, y_pixel, is_in_rays[533]);
assign ray_colors[1067:1066] = GREEN;
square ray_534(534,100 + ((MAX_HEIGHT - 184) / 2),1,184, x_pixel, y_pixel, is_in_rays[534]);
assign ray_colors[1069:1068] = GREEN;
square ray_535(535,100 + ((MAX_HEIGHT - 185) / 2),1,185, x_pixel, y_pixel, is_in_rays[535]);
assign ray_colors[1071:1070] = GREEN;
square ray_536(536,100 + ((MAX_HEIGHT - 186) / 2),1,186, x_pixel, y_pixel, is_in_rays[536]);
assign ray_colors[1073:1072] = GREEN;
square ray_537(537,100 + ((MAX_HEIGHT - 186) / 2),1,186, x_pixel, y_pixel, is_in_rays[537]);
assign ray_colors[1075:1074] = GREEN;
square ray_538(538,100 + ((MAX_HEIGHT - 187) / 2),1,187, x_pixel, y_pixel, is_in_rays[538]);
assign ray_colors[1077:1076] = GREEN;
square ray_539(539,100 + ((MAX_HEIGHT - 188) / 2),1,188, x_pixel, y_pixel, is_in_rays[539]);
assign ray_colors[1079:1078] = GREEN;
square ray_540(540,100 + ((MAX_HEIGHT - 189) / 2),1,189, x_pixel, y_pixel, is_in_rays[540]);
assign ray_colors[1081:1080] = GREEN;
square ray_541(541,100 + ((MAX_HEIGHT - 190) / 2),1,190, x_pixel, y_pixel, is_in_rays[541]);
assign ray_colors[1083:1082] = GREEN;
square ray_542(542,100 + ((MAX_HEIGHT - 191) / 2),1,191, x_pixel, y_pixel, is_in_rays[542]);
assign ray_colors[1085:1084] = GREEN;
square ray_543(543,100 + ((MAX_HEIGHT - 192) / 2),1,192, x_pixel, y_pixel, is_in_rays[543]);
assign ray_colors[1087:1086] = GREEN;
square ray_544(544,100 + ((MAX_HEIGHT - 192) / 2),1,192, x_pixel, y_pixel, is_in_rays[544]);
assign ray_colors[1089:1088] = GREEN;
square ray_545(545,100 + ((MAX_HEIGHT - 193) / 2),1,193, x_pixel, y_pixel, is_in_rays[545]);
assign ray_colors[1091:1090] = GREEN;
square ray_546(546,100 + ((MAX_HEIGHT - 194) / 2),1,194, x_pixel, y_pixel, is_in_rays[546]);
assign ray_colors[1093:1092] = GREEN;
square ray_547(547,100 + ((MAX_HEIGHT - 195) / 2),1,195, x_pixel, y_pixel, is_in_rays[547]);
assign ray_colors[1095:1094] = GREEN;
square ray_548(548,100 + ((MAX_HEIGHT - 196) / 2),1,196, x_pixel, y_pixel, is_in_rays[548]);
assign ray_colors[1097:1096] = GREEN;
square ray_549(549,100 + ((MAX_HEIGHT - 197) / 2),1,197, x_pixel, y_pixel, is_in_rays[549]);
assign ray_colors[1099:1098] = GREEN;
square ray_550(550,100 + ((MAX_HEIGHT - 197) / 2),1,197, x_pixel, y_pixel, is_in_rays[550]);
assign ray_colors[1101:1100] = GREEN;
square ray_551(551,100 + ((MAX_HEIGHT - 198) / 2),1,198, x_pixel, y_pixel, is_in_rays[551]);
assign ray_colors[1103:1102] = GREEN;
square ray_552(552,100 + ((MAX_HEIGHT - 199) / 2),1,199, x_pixel, y_pixel, is_in_rays[552]);
assign ray_colors[1105:1104] = GREEN;
square ray_553(553,100 + ((MAX_HEIGHT - 200) / 2),1,200, x_pixel, y_pixel, is_in_rays[553]);
assign ray_colors[1107:1106] = GREEN;
square ray_554(554,100 + ((MAX_HEIGHT - 201) / 2),1,201, x_pixel, y_pixel, is_in_rays[554]);
assign ray_colors[1109:1108] = GREEN;
square ray_555(555,100 + ((MAX_HEIGHT - 202) / 2),1,202, x_pixel, y_pixel, is_in_rays[555]);
assign ray_colors[1111:1110] = GREEN;
square ray_556(556,100 + ((MAX_HEIGHT - 202) / 2),1,202, x_pixel, y_pixel, is_in_rays[556]);
assign ray_colors[1113:1112] = GREEN;
square ray_557(557,100 + ((MAX_HEIGHT - 203) / 2),1,203, x_pixel, y_pixel, is_in_rays[557]);
assign ray_colors[1115:1114] = GREEN;
square ray_558(558,100 + ((MAX_HEIGHT - 204) / 2),1,204, x_pixel, y_pixel, is_in_rays[558]);
assign ray_colors[1117:1116] = GREEN;
square ray_559(559,100 + ((MAX_HEIGHT - 205) / 2),1,205, x_pixel, y_pixel, is_in_rays[559]);
assign ray_colors[1119:1118] = GREEN;
square ray_560(560,100 + ((MAX_HEIGHT - 206) / 2),1,206, x_pixel, y_pixel, is_in_rays[560]);
assign ray_colors[1121:1120] = GREEN;
square ray_561(561,100 + ((MAX_HEIGHT - 207) / 2),1,207, x_pixel, y_pixel, is_in_rays[561]);
assign ray_colors[1123:1122] = GREEN;
square ray_562(562,100 + ((MAX_HEIGHT - 207) / 2),1,207, x_pixel, y_pixel, is_in_rays[562]);
assign ray_colors[1125:1124] = GREEN;
square ray_563(563,100 + ((MAX_HEIGHT - 208) / 2),1,208, x_pixel, y_pixel, is_in_rays[563]);
assign ray_colors[1127:1126] = GREEN;
square ray_564(564,100 + ((MAX_HEIGHT - 209) / 2),1,209, x_pixel, y_pixel, is_in_rays[564]);
assign ray_colors[1129:1128] = GREEN;
square ray_565(565,100 + ((MAX_HEIGHT - 210) / 2),1,210, x_pixel, y_pixel, is_in_rays[565]);
assign ray_colors[1131:1130] = GREEN;
square ray_566(566,100 + ((MAX_HEIGHT - 211) / 2),1,211, x_pixel, y_pixel, is_in_rays[566]);
assign ray_colors[1133:1132] = GREEN;
square ray_567(567,100 + ((MAX_HEIGHT - 212) / 2),1,212, x_pixel, y_pixel, is_in_rays[567]);
assign ray_colors[1135:1134] = GREEN;
square ray_568(568,100 + ((MAX_HEIGHT - 212) / 2),1,212, x_pixel, y_pixel, is_in_rays[568]);
assign ray_colors[1137:1136] = GREEN;
square ray_569(569,100 + ((MAX_HEIGHT - 213) / 2),1,213, x_pixel, y_pixel, is_in_rays[569]);
assign ray_colors[1139:1138] = GREEN;
square ray_570(570,100 + ((MAX_HEIGHT - 214) / 2),1,214, x_pixel, y_pixel, is_in_rays[570]);
assign ray_colors[1141:1140] = GREEN;
square ray_571(571,100 + ((MAX_HEIGHT - 215) / 2),1,215, x_pixel, y_pixel, is_in_rays[571]);
assign ray_colors[1143:1142] = GREEN;
square ray_572(572,100 + ((MAX_HEIGHT - 216) / 2),1,216, x_pixel, y_pixel, is_in_rays[572]);
assign ray_colors[1145:1144] = GREEN;
square ray_573(573,100 + ((MAX_HEIGHT - 217) / 2),1,217, x_pixel, y_pixel, is_in_rays[573]);
assign ray_colors[1147:1146] = GREEN;
square ray_574(574,100 + ((MAX_HEIGHT - 217) / 2),1,217, x_pixel, y_pixel, is_in_rays[574]);
assign ray_colors[1149:1148] = GREEN;
square ray_575(575,100 + ((MAX_HEIGHT - 218) / 2),1,218, x_pixel, y_pixel, is_in_rays[575]);
assign ray_colors[1151:1150] = GREEN;
square ray_576(576,100 + ((MAX_HEIGHT - 219) / 2),1,219, x_pixel, y_pixel, is_in_rays[576]);
assign ray_colors[1153:1152] = GREEN;
square ray_577(577,100 + ((MAX_HEIGHT - 220) / 2),1,220, x_pixel, y_pixel, is_in_rays[577]);
assign ray_colors[1155:1154] = GREEN;
square ray_578(578,100 + ((MAX_HEIGHT - 221) / 2),1,221, x_pixel, y_pixel, is_in_rays[578]);
assign ray_colors[1157:1156] = GREEN;
square ray_579(579,100 + ((MAX_HEIGHT - 222) / 2),1,222, x_pixel, y_pixel, is_in_rays[579]);
assign ray_colors[1159:1158] = GREEN;
square ray_580(580,100 + ((MAX_HEIGHT - 222) / 2),1,222, x_pixel, y_pixel, is_in_rays[580]);
assign ray_colors[1161:1160] = GREEN;
square ray_581(581,100 + ((MAX_HEIGHT - 223) / 2),1,223, x_pixel, y_pixel, is_in_rays[581]);
assign ray_colors[1163:1162] = GREEN;
square ray_582(582,100 + ((MAX_HEIGHT - 224) / 2),1,224, x_pixel, y_pixel, is_in_rays[582]);
assign ray_colors[1165:1164] = GREEN;
square ray_583(583,100 + ((MAX_HEIGHT - 225) / 2),1,225, x_pixel, y_pixel, is_in_rays[583]);
assign ray_colors[1167:1166] = GREEN;
square ray_584(584,100 + ((MAX_HEIGHT - 226) / 2),1,226, x_pixel, y_pixel, is_in_rays[584]);
assign ray_colors[1169:1168] = GREEN;
square ray_585(585,100 + ((MAX_HEIGHT - 227) / 2),1,227, x_pixel, y_pixel, is_in_rays[585]);
assign ray_colors[1171:1170] = GREEN;
square ray_586(586,100 + ((MAX_HEIGHT - 227) / 2),1,227, x_pixel, y_pixel, is_in_rays[586]);
assign ray_colors[1173:1172] = GREEN;
square ray_587(587,100 + ((MAX_HEIGHT - 228) / 2),1,228, x_pixel, y_pixel, is_in_rays[587]);
assign ray_colors[1175:1174] = GREEN;
square ray_588(588,100 + ((MAX_HEIGHT - 229) / 2),1,229, x_pixel, y_pixel, is_in_rays[588]);
assign ray_colors[1177:1176] = GREEN;
square ray_589(589,100 + ((MAX_HEIGHT - 230) / 2),1,230, x_pixel, y_pixel, is_in_rays[589]);
assign ray_colors[1179:1178] = GREEN;
square ray_590(590,100 + ((MAX_HEIGHT - 231) / 2),1,231, x_pixel, y_pixel, is_in_rays[590]);
assign ray_colors[1181:1180] = GREEN;
square ray_591(591,100 + ((MAX_HEIGHT - 232) / 2),1,232, x_pixel, y_pixel, is_in_rays[591]);
assign ray_colors[1183:1182] = GREEN;
square ray_592(592,100 + ((MAX_HEIGHT - 232) / 2),1,232, x_pixel, y_pixel, is_in_rays[592]);
assign ray_colors[1185:1184] = GREEN;
square ray_593(593,100 + ((MAX_HEIGHT - 233) / 2),1,233, x_pixel, y_pixel, is_in_rays[593]);
assign ray_colors[1187:1186] = GREEN;
square ray_594(594,100 + ((MAX_HEIGHT - 234) / 2),1,234, x_pixel, y_pixel, is_in_rays[594]);
assign ray_colors[1189:1188] = GREEN;
square ray_595(595,100 + ((MAX_HEIGHT - 235) / 2),1,235, x_pixel, y_pixel, is_in_rays[595]);
assign ray_colors[1191:1190] = GREEN;
square ray_596(596,100 + ((MAX_HEIGHT - 236) / 2),1,236, x_pixel, y_pixel, is_in_rays[596]);
assign ray_colors[1193:1192] = GREEN;
square ray_597(597,100 + ((MAX_HEIGHT - 237) / 2),1,237, x_pixel, y_pixel, is_in_rays[597]);
assign ray_colors[1195:1194] = GREEN;
square ray_598(598,100 + ((MAX_HEIGHT - 237) / 2),1,237, x_pixel, y_pixel, is_in_rays[598]);
assign ray_colors[1197:1196] = GREEN;
square ray_599(599,100 + ((MAX_HEIGHT - 238) / 2),1,238, x_pixel, y_pixel, is_in_rays[599]);
assign ray_colors[1199:1198] = GREEN;
square ray_600(600,100 + ((MAX_HEIGHT - 239) / 2),1,239, x_pixel, y_pixel, is_in_rays[600]);
assign ray_colors[1201:1200] = GREEN;
square ray_601(601,100 + ((MAX_HEIGHT - 240) / 2),1,240, x_pixel, y_pixel, is_in_rays[601]);
assign ray_colors[1203:1202] = GREEN;
square ray_602(602,100 + ((MAX_HEIGHT - 241) / 2),1,241, x_pixel, y_pixel, is_in_rays[602]);
assign ray_colors[1205:1204] = GREEN;
square ray_603(603,100 + ((MAX_HEIGHT - 242) / 2),1,242, x_pixel, y_pixel, is_in_rays[603]);
assign ray_colors[1207:1206] = GREEN;
square ray_604(604,100 + ((MAX_HEIGHT - 242) / 2),1,242, x_pixel, y_pixel, is_in_rays[604]);
assign ray_colors[1209:1208] = GREEN;
square ray_605(605,100 + ((MAX_HEIGHT - 243) / 2),1,243, x_pixel, y_pixel, is_in_rays[605]);
assign ray_colors[1211:1210] = GREEN;
square ray_606(606,100 + ((MAX_HEIGHT - 244) / 2),1,244, x_pixel, y_pixel, is_in_rays[606]);
assign ray_colors[1213:1212] = GREEN;
square ray_607(607,100 + ((MAX_HEIGHT - 245) / 2),1,245, x_pixel, y_pixel, is_in_rays[607]);
assign ray_colors[1215:1214] = GREEN;
square ray_608(608,100 + ((MAX_HEIGHT - 246) / 2),1,246, x_pixel, y_pixel, is_in_rays[608]);
assign ray_colors[1217:1216] = GREEN;
square ray_609(609,100 + ((MAX_HEIGHT - 247) / 2),1,247, x_pixel, y_pixel, is_in_rays[609]);
assign ray_colors[1219:1218] = GREEN;
square ray_610(610,100 + ((MAX_HEIGHT - 247) / 2),1,247, x_pixel, y_pixel, is_in_rays[610]);
assign ray_colors[1221:1220] = GREEN;
square ray_611(611,100 + ((MAX_HEIGHT - 248) / 2),1,248, x_pixel, y_pixel, is_in_rays[611]);
assign ray_colors[1223:1222] = GREEN;
square ray_612(612,100 + ((MAX_HEIGHT - 249) / 2),1,249, x_pixel, y_pixel, is_in_rays[612]);
assign ray_colors[1225:1224] = GREEN;
square ray_613(613,100 + ((MAX_HEIGHT - 250) / 2),1,250, x_pixel, y_pixel, is_in_rays[613]);
assign ray_colors[1227:1226] = GREEN;
square ray_614(614,100 + ((MAX_HEIGHT - 251) / 2),1,251, x_pixel, y_pixel, is_in_rays[614]);
assign ray_colors[1229:1228] = GREEN;
square ray_615(615,100 + ((MAX_HEIGHT - 251) / 2),1,251, x_pixel, y_pixel, is_in_rays[615]);
assign ray_colors[1231:1230] = GREEN;
square ray_616(616,100 + ((MAX_HEIGHT - 252) / 2),1,252, x_pixel, y_pixel, is_in_rays[616]);
assign ray_colors[1233:1232] = GREEN;
square ray_617(617,100 + ((MAX_HEIGHT - 253) / 2),1,253, x_pixel, y_pixel, is_in_rays[617]);
assign ray_colors[1235:1234] = GREEN;
square ray_618(618,100 + ((MAX_HEIGHT - 254) / 2),1,254, x_pixel, y_pixel, is_in_rays[618]);
assign ray_colors[1237:1236] = GREEN;
square ray_619(619,100 + ((MAX_HEIGHT - 255) / 2),1,255, x_pixel, y_pixel, is_in_rays[619]);
assign ray_colors[1239:1238] = GREEN;
square ray_620(620,100 + ((MAX_HEIGHT - 256) / 2),1,256, x_pixel, y_pixel, is_in_rays[620]);
assign ray_colors[1241:1240] = GREEN;
square ray_621(621,100 + ((MAX_HEIGHT - 256) / 2),1,256, x_pixel, y_pixel, is_in_rays[621]);
assign ray_colors[1243:1242] = GREEN;
square ray_622(622,100 + ((MAX_HEIGHT - 257) / 2),1,257, x_pixel, y_pixel, is_in_rays[622]);
assign ray_colors[1245:1244] = GREEN;
square ray_623(623,100 + ((MAX_HEIGHT - 258) / 2),1,258, x_pixel, y_pixel, is_in_rays[623]);
assign ray_colors[1247:1246] = GREEN;
square ray_624(624,100 + ((MAX_HEIGHT - 259) / 2),1,259, x_pixel, y_pixel, is_in_rays[624]);
assign ray_colors[1249:1248] = GREEN;
square ray_625(625,100 + ((MAX_HEIGHT - 260) / 2),1,260, x_pixel, y_pixel, is_in_rays[625]);
assign ray_colors[1251:1250] = GREEN;
square ray_626(626,100 + ((MAX_HEIGHT - 261) / 2),1,261, x_pixel, y_pixel, is_in_rays[626]);
assign ray_colors[1253:1252] = GREEN;
square ray_627(627,100 + ((MAX_HEIGHT - 261) / 2),1,261, x_pixel, y_pixel, is_in_rays[627]);
assign ray_colors[1255:1254] = GREEN;
square ray_628(628,100 + ((MAX_HEIGHT - 262) / 2),1,262, x_pixel, y_pixel, is_in_rays[628]);
assign ray_colors[1257:1256] = GREEN;
square ray_629(629,100 + ((MAX_HEIGHT - 263) / 2),1,263, x_pixel, y_pixel, is_in_rays[629]);
assign ray_colors[1259:1258] = GREEN;
square ray_630(630,100 + ((MAX_HEIGHT - 264) / 2),1,264, x_pixel, y_pixel, is_in_rays[630]);
assign ray_colors[1261:1260] = GREEN;
square ray_631(631,100 + ((MAX_HEIGHT - 265) / 2),1,265, x_pixel, y_pixel, is_in_rays[631]);
assign ray_colors[1263:1262] = GREEN;
square ray_632(632,100 + ((MAX_HEIGHT - 265) / 2),1,265, x_pixel, y_pixel, is_in_rays[632]);
assign ray_colors[1265:1264] = GREEN;
square ray_633(633,100 + ((MAX_HEIGHT - 266) / 2),1,266, x_pixel, y_pixel, is_in_rays[633]);
assign ray_colors[1267:1266] = GREEN;
square ray_634(634,100 + ((MAX_HEIGHT - 267) / 2),1,267, x_pixel, y_pixel, is_in_rays[634]);
assign ray_colors[1269:1268] = GREEN;
square ray_635(635,100 + ((MAX_HEIGHT - 268) / 2),1,268, x_pixel, y_pixel, is_in_rays[635]);
assign ray_colors[1271:1270] = GREEN;
square ray_636(636,100 + ((MAX_HEIGHT - 269) / 2),1,269, x_pixel, y_pixel, is_in_rays[636]);
assign ray_colors[1273:1272] = GREEN;
square ray_637(637,100 + ((MAX_HEIGHT - 269) / 2),1,269, x_pixel, y_pixel, is_in_rays[637]);
assign ray_colors[1275:1274] = GREEN;
square ray_638(638,100 + ((MAX_HEIGHT - 270) / 2),1,270, x_pixel, y_pixel, is_in_rays[638]);
assign ray_colors[1277:1276] = GREEN;
square ray_639(639,100 + ((MAX_HEIGHT - 271) / 2),1,271, x_pixel, y_pixel, is_in_rays[639]);
assign ray_colors[1279:1278] = GREEN;

endmodule

